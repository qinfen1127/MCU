//==========================================================================================================================
//  @File Name  :  temp.v
//  @File Type  :  verilog
//  @Author     :  Howard
//  @E-mail     :  qinfen1127@163.com
//  @Date       :  2024-07-06
//  @Function   :  just make a test
//==========================================================================================================================

module temp #(

)(

);


endmodule

